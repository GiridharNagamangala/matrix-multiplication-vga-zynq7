`timescale 1ns / 1ps
module vga_digit_rom (
    input        clk,
    input  [3:0] digit_code, // 0–9
    input  [3:0] row,        // 0–15
    input  [2:0] col,        // 0–7
    output wire  pixel
);

    reg [7:0] rom [0:12][0:15];

    always @(posedge clk) begin
        // Zero
        rom [0][0] <= 8'h00; rom [0][1] <= 8'h00; rom [0][2] <= 8'h7c; rom [0][3] <= 8'h66;
        rom [0][4] <= 8'h66; rom [0][5] <= 8'h66; rom [0][6] <= 8'h66; rom [0][7] <= 8'h66;
        rom [0][8] <= 8'h66; rom [0][9] <= 8'h66; rom [0][10] <= 8'h66; rom [0][11] <= 8'h66;
        rom [0][12] <= 8'h7c; rom [0][13] <= 8'h00; rom [0][14] <= 8'h00; rom [0][15] <= 8'h00;

        //One
        rom [1][0] <= 8'h00; rom [1][1] <= 8'h00; rom [1][2] <= 8'h18; rom [1][3] <= 8'h38;
        rom [1][4] <= 8'h18; rom [1][5] <= 8'h18; rom [1][6] <= 8'h18; rom [1][7] <= 8'h18;
        rom [1][8] <= 8'h18; rom [1][9] <= 8'h18; rom [1][10] <= 8'h18; rom [1][11] <= 8'h18;
        rom [1][12] <= 8'h7e; rom [1][13] <= 8'h00; rom [1][14] <= 8'h00; rom [1][15] <= 8'h00;

        // Two
        rom [2][0] <= 8'h00; rom [2][1] <= 8'h00; rom [2][2] <= 8'h7c; rom [2][3] <= 8'h66;
        rom [2][4] <= 8'h60; rom [2][5] <= 8'h30; rom [2][6] <= 8'h18; rom [2][7] <= 8'h0c;
        rom [2][8] <= 8'h0c; rom [2][9] <= 8'h66; rom [2][10] <= 8'h66; rom [2][11] <= 8'h66;
        rom [2][12] <= 8'h7c; rom [2][13] <= 8'h00; rom [2][14] <= 8'h00; rom [2][15] <= 8'h00;

        // Three
        rom [3][0] <= 8'h00; rom [3][1] <= 8'h00; rom [3][2] <= 8'h7c; rom [3][3] <= 8'h66;
        rom [3][4] <= 8'h06; rom [3][5] <= 8'h3c; rom [3][6] <= 8'h06; rom [3][7] <= 8'h06;
        rom [3][8] <= 8'h66; rom [3][9] <= 8'h66; rom [3][10] <= 8'h66; rom [3][11] <= 8'h66;
        rom [3][12] <= 8'h7c; rom [3][13] <= 8'h00; rom [3][14] <= 8'h00; rom [3][15] <= 8'h00;

        // Four
        rom [4][0] <= 8'h00; rom [4][1] <= 8'h00; rom [4][2] <= 8'h18; rom [4][3] <= 8'h38;
        rom [4][4] <= 8'h68; rom [4][5] <= 8'h38; rom [4][6] <= 8'hfe; rom [4][7] <= 8'h08;
        rom [4][8] <= 8'h08; rom [4][9] <= 8'h08; rom [4][10] <= 8'h08; rom [4][11] <= 8'h08;
        rom [4][12] <= 8'hfe; rom [4][13] <= 8'h00; rom [4][14] <= 8'h00; rom [4][15] <= 8'h00;

        // Five
        rom [5][0] <= 8'h00; rom [5][1] <= 8'h00; rom [5][2] <= 8'hfc; rom [5][3] <= 8'hc0;
        rom [5][4] <= 8'hc0; rom [5][5] <= 8'hc0; rom [5][6] <= 8'hf8; rom [5][7] <= 8'h06;
        rom [5][8] <= 8'h06; rom [5][9] <= 8'h06; rom [5][10] <= 8'h66; rom [5][11] <= 8'h66;
        rom [5][12] <= 8'h7c; rom [5][13] <= 8'h00; rom [5][14] <= 8'h00; rom [5][15] <= 8'h00;

        // Six
        rom [6][0] <= 8'h00; rom [6][1] <= 8'h00; rom [6][2] <= 8'h7c; rom [6][3] <= 8'h66;
        rom [6][4] <= 8'h60; rom [6][5] <= 8'hc0; rom [6][6] <= 8'hf8; rom [6][7] <= 8'h66;
        rom [6][8] <= 8'h66; rom [6][9] <= 8'h66; rom [6][10] <= 8'h66; rom [6][11] <= 8'h66;
        rom [6][12] <= 8'h7c; rom [6][13] <= 8'h00; rom [6][14] <= 8'h00; rom [6][15] <= 8'h00;

        // Seven
        rom [7][0] <= 8'h00; rom [7][1] <= 8'h00; rom [7][2] <= 8'hfe; rom [7][3] <= 8'h66;
        rom [7][4] <= 8'h06; rom [7][5] <= 8'h0c; rom [7][6] <= 8'h18; rom [7][7] <= 8'h30;
        rom [7][8] <= 8'h60; rom [7][9] <= 8'h60; rom [7][10] <= 8'h60; rom [7][11] <= 8'h60;
        rom [7][12] <= 8'h60; rom [7][13] <= 8'h00; rom [7][14] <= 8'h00; rom [7][15] <= 8'h00;

        // Eight
        rom [8][0] <= 8'h00; rom [8][1] <= 8'h00; rom [8][2] <= 8'h7c; rom [8][3] <= 8'h66;
        rom [8][4] <= 8'h66; rom [8][5] <= 8'h66; rom [8][6] <= 8'h7c; rom [8][7] <= 8'h66;
        rom [8][8] <= 8'h66; rom [8][9] <= 8'h66; rom [8][10] <= 8'h66; rom [8][11] <= 8'h66;
        rom [8][12] <= 8'h7c; rom [8][13] <= 8'h00; rom [8][14] <= 8'h00; rom [8][15] <= 8'h00;

        // Nine
        rom [9][0] <= 8'h00; rom [9][1] <= 8'h00; rom [9][2] <= 8'h7c; rom [9][3] <= 8'h66;
        rom [9][4] <= 8'h66; rom [9][5] <= 8'h66; rom [9][6] <= 8'h7c; rom [9][7] <= 8'h06;
        rom [9][8] <= 8'h06; rom [9][9] <= 8'h06; rom [9][10] <= 8'h06; rom [9][11] <= 8'h06;
        rom [9][12] <= 8'h7c; rom [9][13] <= 8'h00; rom [9][14] <= 8'h00; rom [9][15] <= 8'h00;

        // multiplication symbol
        rom [10][0] <= 8'h00; rom [10][1] <= 8'h00; rom [10][2] <= 8'h00; rom [10][3] <= 8'h00;
        rom [10][4] <= 8'h81; rom [10][5] <= 8'h42; rom [10][6] <= 8'h24; rom [10][7] <= 8'h18;
        rom [10][8] <= 8'h18; rom [10][9] <= 8'h24; rom [10][10] <= 8'h42; rom [10][11] <= 8'h81;
        rom [10][12] <= 8'h00; rom [10][13] <= 8'h00; rom [10][14] <= 8'h00; rom [10][15] <= 8'h00;

        // Equals symbol
        rom [11][0] <= 8'h00; rom [11][1] <= 8'h00; rom [11][2] <= 8'h00; rom [11][3] <= 8'h00;
        rom [11][4] <= 8'h00; rom [11][5] <= 8'hff; rom [11][6] <= 8'hff; rom [11][7] <= 8'h00;
        rom [11][8] <= 8'h00; rom [11][9] <= 8'hff; rom [11][10] <= 8'hff; rom [11][11] <= 8'h00;
        rom [11][12] <= 8'h00; rom [11][13] <= 8'h00; rom [11][14] <= 8'h00; rom [11][15] <= 8'h00;

        // Decimal point
        rom [12][0] <= 8'h00; rom [12][1] <= 8'h00; rom [12][2] <= 8'h00; rom [12][3] <= 8'h00;
        rom [12][4] <= 8'h00; rom [12][5] <= 8'h00; rom [12][6] <= 8'h00; rom [12][7] <= 8'h00;
        rom [12][8] <= 8'h00; rom [12][9] <= 8'h00; rom [12][10] <= 8'h00; rom [12][11] <= 8'h18;
        rom [12][12] <= 8'h18; rom [12][13] <= 8'h00; rom [12][14] <= 8'h00; rom [12][15] <= 8'h00;

    end

    assign pixel = rom[digit_code][row][col];

endmodule
